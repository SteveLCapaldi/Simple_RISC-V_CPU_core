`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/05/07 19:54:24
// Design Name: 
// Module Name: rom1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rom1 #(  
    parameter DWIDTH = 32,  
    parameter AWIDTH = 32,  
    parameter DEPTH  = 32  
)(  
    input rst,  
    input [AWIDTH - 1 : 0] PC,  
    input en_fetch,  
    output reg [DWIDTH - 1 : 0] instruction
    //output reg en_in  
);  
    reg [DWIDTH - 1 : 0] mem[0 : DEPTH - 1];  
  
    initial begin  
        // ��ʼ��ROM���ݣ���ʾ����  
       /* mem[0] = 32'h0000_0000; //inst=0 
        mem[1] = 32'h0000_0037; // LUI,��r0��Ϊ��ַ�Ĵ������һ�ַΪ0
        mem[2] = 32'h0000_2083;//LW,����ڴ��ַ0������λ���ϵ�ֵ����r1(r1=1)
        mem[3] = 32'h0000_A103;//LW,����ڴ��ַ1������λ���ϵ�ֵ����r2(r2=2)
        mem[4] = 32'h0001_2183;//LW,����ڴ��ַ2������λ���ϵ�ֵ����r3(r3=3)
        mem[5] = 32'h0012_1163;//BNE,ƫ����Ϊ2��
        mem[6] = 32'h0010_8093;//ADDI,r1�ټ���1��r1=2)
        mem[7] = 32'h0010_8113;//ADDI,r1�ټ���1��r2(r2=3) 
        mem[8] = 32'h0020_D083;//ADD,r1����r2���ٸ�r1(r1=5)     
        // ... ������ַ�ĳ�ʼ��  */
        mem[0] = 32'h0000_0000; //inst=0
        mem[1] = 32'b00000000000000000000000000110111;//  LUI 0
        mem[2] = 32'b00000000000100000010000010000011;//LW��1load���Ĵ�����ַ1 000000000001  00000 010 00001 0000011
        mem[3] = 32'b00000000001000000010000100000011;//LW��2load��Ĵ�����ַ2 000000000010  00000 010 00010 0000011
        mem[4] = 32'b0000000_00001_00001_010_00011_0100011;//SW���Ĵ���1��ֵ����Ĵ���1�ĵ�ַ+2��ram 0000000 00001 00001 010 00011 0100011
       // mem[4] = 32'b00000000000100001000000010010011;//addi �Ĵ���1��ֵ��������1��Ӳ����ڼĴ���1 32'b000000000001 00001 000 00001 0010011
        //mem[5] = 32'b00000000001000001000000110110011 ;//ADD���Ĵ���1�ӼĴ���2���ڼĴ���3 32'b0000000 00010 00001 000 00011 0110011 
       // mem[6] = 32'b01000000000100011000001000110011 ;//SUB�Ĵ���3���Ĵ���1�����ڼĴ���4 32'b 0100000 00011 00001 000 00100 0110011 
        //mem[7] = 32'b0_0_000000_00011_00100_000_0010_0_1100011;//BEQ���Ĵ���3�ͼĴ���4�Ƚ�offset��2
        //mem[7] = 32'b0_0_000000_00011_00100_001_0001_0_1100011;//BNE���Ĵ���3�ͼĴ���4�Ƚ�offset��2
        //mem[7] = 32'b000000000010_00001_000_01001_1100111;//JALR �Ĵ���1��ֵ����PC��Ϊ��PC����PC+1����Ĵ���9
       // mem[7] = 32'b0_0000000010_0_00000000_01001_1101111;//JAL PC+immm(2)��pc+1����Ĵ���9
        //mem[7]= 32'b0000000_00001_00010_001_01001_0110011;//SLL���Ĵ���2���ƼĴ���1��2λ�����ڼĴ���9
        //mem[7] = 32'b0000000_00010_00001_001_01010_0010011;//SLLI,�Ĵ���1����2λ�����ڼĴ���10
        
       // mem[8] = 32'b0000000_00011_00001_010_00101_0110011;// SLT���Ĵ���1�ͼĴ���3�Ƚϣ��Ĵ���5��һ
       // mem[9] = 32'b0000000_00001_00011_010_00110_0110011;// SLT���Ĵ���3�ͼĴ���1�Ƚϣ��Ĵ���6��0
        //mem[10] = 32'b000000000111_00001_111_00111_0010011;//ANDI �Ĵ���1��������7�룬���ڼĴ���7
        //mem[11] = 32'b000000011000_00001_100_01000_0010011;//XORI �Ĵ���1��������24��򣬴��ڼĴ���8
        //mem[12] = 32'b000000000010_00001_000_01001_1100111;//JALR �Ĵ���1��ֵ����PC��Ϊ��PC����PC+1����Ĵ���9
    end  

    always @(*) begin  
        if (rst == 1) begin  
            // ��λʱ�������Чָ���validΪ0  
            instruction = 0;  
        end else if (en_fetch) begin  
            // ���readyΪ�� 
            instruction = mem[PC];

        end else begin  
            // ���readyΪ�ͣ�����ȡ��ָ��
            // ���ﲻ��Ҫ���κ����飬��Ϊinstruction��valid��rst��readyΪ����������Ѿ���������  
        end  
    end  
  
endmodule